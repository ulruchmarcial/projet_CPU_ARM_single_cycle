-- instruction_memory.vhd
library ieee;
use ieee.std_logic_1164.all;
--use ieee.numeric_std_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity instruction_memory is
  port (
    A : in  std_logic_vector(4 downto 0);  -- PC(6 downto 2)
    RD : out std_logic_vector(31 downto 0)  -- instruction lues
  );
end entity;

architecture rtl of instruction_memory is
  type mem_type is array (0 to 31) of std_logic_vector(31 downto 0);
  signal rom : mem_type := (
    0 => "11100000010000000000000000000000",  -- SUB r0, r0, r0 
    1 => "11100010100000000101000000001000",   -- ADD r5,r0, #8
    2 => "11100010010001010011000000000011",   -- SUB r3,r5, #3
    3 => "11100001010100110000000000000101",   -- CMP r3, r5 
    4 => "11100001101000000100000100000011",   -- MOV r4, r3, LSL #2
    5 => "11100011010101000110000000001100",   -- CMP R4, #12
    6 => "11100010100000110110000000011110",   -- ADD R6, R3, #30
    7 => "11100001101000000000001110000110",   -- LSL R0, R6, #7
    8 => "11100101100100110111000000000100",   -- LDR R7, [R3, #8]
    9 => "11100001101000001000101011100101",   -- ROR R8, R5, #21
   --10 => "11100001101000001000101011100101",   -- ROR R8, R5, #21
    --11 => "10110010100001010111000000000001",   --ADDLT r7, r5, #1 
    --12 => "11100000010001110111000000000010",   --  AND r7, r7, r2
    --13 => "11100101100000110111000001010100",   --STR r7, [r3, #84]
    --14 => "11100101100100000010000001100000",   --STR r2, [r0, #96]
    --15 => "11100000100010000101000000000000",   --ADD r5, r8, #0 
    --16 => "11100010100000000010000000001110",   --MOV r2, #14 
    --17 => "11100010100000000010000000001101",   --MOV r2, #13
    --18 => "11100010100000000010000000001010",   -- MOV r2, #10
    --19 => "11100101100000000010000001100100",   -- STR r2, [r0, #100] 
   -- Instructions suppl�mentaires pour tester CMP, LSL, LSR, ASR, ROR
    --20 => "11100010100000000110000000001000", -- MOV r6, #8
   -- 21 => "11100001010100100000000000000110", -- CMP r2, r6
   -- 22 => "11001010100000001001000000000001", -- MOVGT r9, #1
   -- 23 => "11010010100000001001000000000000", -- MOVLE r9, #0
   -- 24 => "11100010100000000001000000010000", -- MOV r1, #16
   -- 25 => "11100001101000001010000100000001", -- LSL r10, r1, #2
   -- 26 => "11100001101000001011000100100001", -- LSR r11, r1, #2
   -- 27 => "11100010100000001100000011110000", -- MOV r12, #240
   -- 28 => "11100001101000001101001001000000", -- ASR r13, r12, #4 (r13 = 240 >> 4 = 15)
    --29 => "11100001101000001110000101100000", -- ROR r14, r12, #4 (rotation droite)
    --30 => "11100001010101010000000000001011", -- CMP r10, r11
   -- 31 => "00000010100000001111000001100011", -- MOVEQ r15, #99
    --32 => "11100001101000100100001100010010", -- LSL r4, r2, r3
   -- 33 => "11100001101000100101001100110010", -- LSR r5, r2, r3
    --34 => "11100001101000100110001101010010", -- ASR r6, r2, r3
   -- 35 => "11100001101000100111001101110010", -- ROR r7, r2, r3
   -- 36 => "11100011010101110000000000000000", -- CMP r7, #0
   -- 37 => "00010010100010001000000000000001", -- ADDNE r8, r8, #1
    --38 => "11100101100000001010000001101000", -- STR r10, [r0, #104]
   -- 39 => "11100101100000001110000001101100", -- STR r14, [r0, #108]
    others => (others => '0')
  );
begin
  RD <= rom(to_integer(unsigned(A)));
end architecture;
